module vending_machine (
    input  logic clk,
    input  logic rst_n,    // Active low reset
    input  logic nickel,   // 5 cents
    input  logic dime,     // 10 cents
    output logic dispense, // Merchandise out
    output logic change    // 5 cent nickel change
);

    // TODO: Implement the vending machine logic here

endmodule